module disp(
    Clk,
    Reset_n,
    Disp_Data,
    SEL,
    SEG
);
    input Clk;
    input Reset_n;
    input [7:0] Disp_Data; // 8 bits for 2 digits
    output reg [1:0] SEL;   // Only 2 digits
    output reg [7:0] SEG;
    
    parameter MCNT_1MS = 1000000 /20 - 1;
    parameter MCNT_SEL = 2 - 1; // 2 digits
    reg [15:0] cnt_1ms;
    reg [1:0] cnt_sel; // Change to 2-bit counter for 2 digits
    reg [1:0] encode_sel;
    reg [7:0] LUT_seg;
    reg [3:0] data_temp;

    // 1ms Counter
    always @(posedge Clk or negedge Reset_n) begin
        if (!Reset_n)
            cnt_1ms <= 0;
        else if (cnt_1ms == MCNT_1MS)
            cnt_1ms <= 0;
        else 
            cnt_1ms <= cnt_1ms + 1'b1;
    end

    // Digit Selection Counter
    always @(posedge Clk or negedge Reset_n) begin
        if (!Reset_n)
            cnt_sel <= 0;
        else if (cnt_1ms == MCNT_1MS) begin
            if (cnt_sel == MCNT_SEL)
                cnt_sel <= 0;
            else
                cnt_sel <= cnt_sel + 1'b1;
        end
    end

    // 2-to-4 Decoder
    always @(*) begin
        case (cnt_sel)
            2'b00: encode_sel = 2'b01; // Select first digit
            2'b01: encode_sel = 2'b10; // Select second digit
        endcase
    end

    always @(posedge Clk or negedge Reset_n) begin
        if (!Reset_n)
            SEL <= 0;
        else
            SEL <= encode_sel;
    end

    // Segment Selection
    always @(*) begin
        case (cnt_sel)
            2'b00: data_temp = Disp_Data[3:0]; // First digit
            2'b01: data_temp = Disp_Data[7:4]; // Second digit
        endcase
    end

    // Segment Encoding
    always @(*) begin
        case (data_temp)
            0  : LUT_seg = 8'hc0; // 0
            1  : LUT_seg = 8'hf9; // 1
            2  : LUT_seg = 8'ha4; // 2
            3  : LUT_seg = 8'hb0; // 3
            4  : LUT_seg = 8'h99; // 4
            5  : LUT_seg = 8'h92; // 5
            6  : LUT_seg = 8'h82; // 6
            7  : LUT_seg = 8'hf8; // 7
            8  : LUT_seg = 8'h80; // 8
            9  : LUT_seg = 8'h90; // 9
            4'ha: LUT_seg = 8'h88; // A
            4'hb: LUT_seg = 8'h83; // b
            4'hc: LUT_seg = 8'hc6; // C
            4'hd: LUT_seg = 8'ha1; // d
            4'he: LUT_seg = 8'h86; // E
            4'hf: LUT_seg = 8'h8e; // F
            default: LUT_seg = 8'hff; // Off
        endcase
    end

    always @(posedge Clk or negedge Reset_n) begin
        if (!Reset_n)
            SEG <= 0;
        else
            SEG <= LUT_seg;  
    end

endmodule